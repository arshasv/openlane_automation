module top;
initial begin
    $display("Hello, Verilog!");
    $finish;
end
endmodule
